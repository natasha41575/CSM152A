module 4_bit_counter ();

// Declaring registers for 4 D Flip-Flops
reg reg_1;